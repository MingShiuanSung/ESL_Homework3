`timescale 1ps / 1ps
/*****************************************************************************
    Verilog RTL Description
    
    Configured at: 14:46:16 CST (+0800), Tuesday 12 April 2022
    Configured on: ws37
    Configured by: u107061139 (u107061139)
    
    Created by: Stratus DpOpt 2019.1.01 
*******************************************************************************/

module GaussFilter_N_Mux_2_2_2_4 (
	ctrl1,
	out1
	); /* architecture "behavioural" */ 
input  ctrl1;
output [1:0] out1;
wire [1:0] asc001;

reg [1:0] asc001_tmp_0;
assign asc001 = asc001_tmp_0;
always @ (ctrl1) begin
	case (ctrl1)
		1'B1 : asc001_tmp_0 = 2'B11 ;
		default : asc001_tmp_0 = 2'B00 ;
	endcase
end

assign out1 = asc001;
endmodule

/* CADENCE  uLD5Twk= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE ******/


